library verilog;
use verilog.vl_types.all;
entity JSQ_FZN_top_vlg_vec_tst is
end JSQ_FZN_top_vlg_vec_tst;
