module part4_demo( 
	input [7:0] add_sub,
	input [7:0] dataa,
	input [7:0] datab,
	output overflow,
	output [7:0] result);
part4_add demo(
	add_sub,
	dataa,
	datab,
	overflow,
	result);
endmodule 
	