module ls47(input [15:0]sw,output [6:0] hex3,
                output [6:0] hex2,hex1,hex0); 
					 
//实际上，此程序还有修正空间，逻辑与可以用乘法代替，逻辑或可以用加法，能缩减程序长度
//工作原理与74ls47类似，需要改变的是1010-1111时gfedcba=1111111,即全灭					 
assign hex0[0]=( (~sw[3])&(~sw[2])&(~sw[1])&sw[0] )|( sw[3]&sw[1] )| ( sw[2]&(~sw[0]))|(sw[3]*sw[2]+sw[3]*sw[1]);
assign hex0[1]=( sw[3]&sw[1]) | ( sw[2]&sw[1]&(~sw[0])) | ( sw[2]&sw[0]&(~sw[1]))|(sw[3]*sw[2]+sw[3]*sw[1]);
assign hex0[2]=( sw[3]&sw[2]) | ( sw[1]&(~sw[2])&(~sw[0]))|(sw[3]*sw[2]+sw[3]*sw[1]);
assign hex0[3]=( sw[2]&sw[1]&sw[0]) |( sw[2]&(~sw[1])&(~sw[0])) |( sw[0]&(~sw[2])&(~sw[1]))|(sw[3]*sw[2]+sw[3]*sw[1]);
assign hex0[4]=( sw[2]&(~sw[1])) | sw[0]|(sw[3]*sw[2]+sw[3]*sw[1]);
assign hex0[5]=( (~sw[3])&(~sw[2])&sw[0]) |( (~sw[2]&sw[1])) |( sw[1]&sw[0])|(sw[3]*sw[2]+sw[3]*sw[1]);
assign hex0[6]=( (~sw[3])&(~sw[2])&(~sw[1])) |( sw[2]&sw[1]&sw[0])|(sw[3]*sw[2]+sw[3]*sw[1]);
//再处理其他数码管，逻辑上类似，加4即可
assign hex1[0]=( (~sw[3+4])&(~sw[2+4])&(~sw[1+4])&sw[0+4] )|( sw[3+4]&sw[1+4] )| ( sw[2+4]&(~sw[0+4]))|(sw[3+4]*sw[2+4]+sw[3+4]*sw[1+4]);
assign hex1[1]=( sw[3+4]&sw[1+4]) | ( sw[2+4]&sw[1+4]*(~sw[0+4])) | ( sw[2+4]&sw[0+4]&(~sw[1+4]))|(sw[3+4]*sw[2+4]+sw[3+4]*sw[1+4]);
assign hex1[2]=( sw[3+4]&sw[2+4]) | ( sw[1+4]&(~sw[2+4])&(~sw[0+4]))|(sw[3+4]*sw[2+4]+sw[3+4]*sw[1+4]);
assign hex1[3]=( sw[2+4]&sw[1+4]&sw[0+4]) |( sw[2+4]&(~sw[1+4])&(~sw[0+4])) |( sw[0+4]&(~sw[2+4])&(~sw[1+4]))|(sw[3+4]*sw[2+4]+sw[3+4]*sw[1+4]);
assign hex1[4]=( sw[2+4]&(~sw[1+4])) | sw[0+4]|(sw[3+4]*sw[2+4]+sw[3+4]*sw[1+4]);
assign hex1[5]=( (~sw[3+4])&(~sw[2+4])&sw[0+4]) |( (~sw[2+4]&sw[1+4])) |( sw[1+4]&sw[0+4])|(sw[3+4]*sw[2+4]+sw[3+4]*sw[1+4]);
assign hex1[6]=( (~sw[3+4])&(~sw[2+4])&(~sw[1+4])) |( sw[2+4]&sw[1+4]&sw[0+4])|(sw[3+4]*sw[2+4]+sw[3+4]*sw[1+4]);
//再加4
assign hex2[0]=( (~sw[3+8])&(~sw[2+8])&(~sw[1+8])&sw[0+8] )|( sw[3+8]&sw[1+8] )| ( sw[2+8]&(~sw[0+8]))|(sw[3+8]*sw[2+8]+sw[3+8]*sw[1+8]);
assign hex2[1]=( sw[3+8]&sw[1+8]) | ( sw[2+8]&sw[1+8]*(~sw[0+8])) | ( sw[2+8]&sw[0+8]&(~sw[1+8]))|(sw[3+8]*sw[2+8]+sw[3+8]*sw[1+8]);
assign hex2[2]=( sw[3+8]&sw[2+8]) | ( sw[1+8]&(~sw[2+8])&(~sw[0+8]))|(sw[3+8]*sw[2+8]+sw[3+8]*sw[1+8]);
assign hex2[3]=( sw[2+8]&sw[1+8]&sw[0+8]) |( sw[2+8]&(~sw[1+8])&(~sw[0+8])) |( sw[0+8]&(~sw[2+8])&(~sw[1+8]))|(sw[3+8]*sw[2+8]+sw[3+8]*sw[1+8]);
assign hex2[4]=( sw[2]&(~sw[1])) | sw[0]|(sw[3+8]*sw[2+8]+sw[3+8]*sw[1+8]);
assign hex2[5]=( (~sw[3+8])&(~sw[2+8])&sw[0+8]) |( (~sw[2+8]&sw[1+8])) |( sw[1+8]&sw[0+8])|(sw[3+8]*sw[2+8]+sw[3+8]*sw[1+8]);
assign hex2[6]=( (~sw[3+8])&(~sw[2+8])&(~sw[1+8])) |( sw[2+8]&sw[1+8]&sw[0+8])|(sw[3+8]*sw[2+8]+sw[3+8]*sw[1+8]);
//加4
assign hex3[0]=( (~sw[3+12])&(~sw[2+12])&(~sw[1+12])&sw[0+12] )|( sw[3+12]&sw[1+12] )| ( sw[2+12]&(~sw[0+12]))|(sw[3+12]*sw[2+12]+sw[3+12]*sw[1+12]);
assign hex3[1]=( sw[3+12]&sw[1+12]) | ( sw[2+12]&sw[1+12]*(~sw[0+12])) | ( sw[2+12]&sw[0+12]&(~sw[1+12]))|(sw[3+12]*sw[2+12]+sw[3+12]*sw[1+12]);
assign hex3[2]=( sw[3+12]&sw[2+12]) | ( sw[1+12]&(~sw[2+12])&(~sw[0+12]))|(sw[3+12]*sw[2+12]+sw[3+12]*sw[1+12]);
assign hex3[3]=( sw[2+12]&sw[1+12]&sw[0+12]) |( sw[2+12]&(~sw[1+12])&(~sw[0+12])) |( sw[0+12]&(~sw[2+12])&(~sw[1+12]))|(sw[3+12]*sw[2+12]+sw[3+12]*sw[1+12]);
assign hex3[4]=( sw[2+12]&(~sw[1+12])) | sw[0+12]|(sw[3+12]*sw[2+12]+sw[3+12]*sw[1+12]);
assign hex3[5]=( (~sw[3+12])&(~sw[2+12])&sw[0+12]) |( (~sw[2+12]&sw[1])) |( sw[1+12]&sw[0+12])|(sw[3+12]*sw[2+12]+sw[3+12]*sw[1+12]);
assign hex3[6]=( (~sw[3+12])&(~sw[2+12])&(~sw[1+12])) |( sw[2+12]&sw[1+12]&sw[0+12])|(sw[3+12]*sw[2+12]+sw[3+12]*sw[1+12]);
endmodule 
