library verilog;
use verilog.vl_types.all;
entity lab3_part3_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        d               : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end lab3_part3_vlg_sample_tst;
